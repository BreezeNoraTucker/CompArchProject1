`timescale 1ns / 1ns
`include "FlowControl.v"

module LDC (input [63:0][19:0] mem, input C, input[5:0] R, output wire [19:0] out);    
    MUX()
endmodule