`timescale 1ns / 1ns
`include "FlowControl.v"

// MUX TESTBENCH
module MUX_tb;

reg [31:0][19:0] a;
reg [4:0] sel;
wire [19:0] out;


MUX multi(a,sel,out);

initial begin

    $dumpfile("FlowControl.vcd");
    $dumpvars(0, MUX_tb);
    a[0] = 20'b00000000000000000000;
    a[1] = 20'b00000000000000000001;
    a[2] = 20'b00000000000000000010;
    a[3] = 20'b00000000000000000011;
    a[4] = 20'b00000000000000000100;
    a[5] = 20'b00000000000000000101;
    a[6] = 20'b00000000000000000110;
    a[7] = 20'b00000000000000000111;
    a[8] = 20'b00000000000000001000;
    a[9] = 20'b00000000000000001001;
    a[10] = 20'b00000000000000001010;
    a[11] = 20'b00000000000000001011;
    a[12] = 20'b00000000000000001100;
    a[13] = 20'b00000000000000001101;
    a[14] = 20'b00000000000000001110;
    a[15] = 20'b00000000000000001111;
    a[16] = 20'b00000000000000010000;
    a[17] = 20'b00000000000000010001;
    a[18] = 20'b00000000000000010010;
    a[19] = 20'b00000000000000010011;
    a[20] = 20'b00000000000000010100;
    a[21] = 20'b00000000000000010101;
    a[22] = 20'b00000000000000010110;
    a[23] = 20'b00000000000000010111;
    a[24] = 20'b00000000000000011000;
    a[25] = 20'b00000000000000011001;
    a[26] = 20'b00000000000000011010;
    a[27] = 20'b00000000000000011011;
    a[28] = 20'b00000000000000011100;
    a[29] = 20'b00000000000000011101;
    a[30] = 20'b00000000000000011110;
    a[31] = 20'b00000000000000011111;

    sel = 5'b00000;
    #10;

    sel = 5'b00001;
    #10;
    
    sel = 5'b00010;
    #10;

    sel = 5'b00100;
    #10;

    sel = 5'b11111;
    #10;

    $display("test complete");
    $finish;

end

endmodule