`timescale 1ns / 1ns
`include "../MemoryBank.v"

// MEMORY BANK LOADING CONSTANT TESTBENCH
module LDC_tb;

reg [63:0][19:0] a;
reg [19:0] C;
reg [5:0] R;
wire [19:0] out;
wire [19:0] buff1;
wire [19:0] buff2;


LDC mem(a,C,R,out,buff1,buff2);

initial begin

    $dumpfile("MemoryBank.vcd");
    $dumpvars(0, LDC_tb);
    a[0] = 20'b00000000000000000000;
    a[1] = 20'b00000000000000000001;
    a[2] = 20'b00000000000000000010;
    a[3] = 20'b00000000000000000011;
    a[4] = 20'b00000000000000000100;
    a[5] = 20'b00000000000000000101;
    a[6] = 20'b00000000000000000110;
    a[7] = 20'b00000000000000000111;
    a[8] = 20'b00000000000000001000;
    a[9] = 20'b00000000000000001001;
    a[10] = 20'b00000000000000001010;
    a[11] = 20'b00000000000000001011;
    a[12] = 20'b00000000000000001100;
    a[13] = 20'b00000000000000001101;
    a[14] = 20'b00000000000000001110;
    a[15] = 20'b00000000000000001111;
    a[16] = 20'b00000000000000010000;
    a[17] = 20'b00000000000000010001;
    a[18] = 20'b00000000000000010010;
    a[19] = 20'b00000000000000010011;
    a[20] = 20'b00000000000000010100;
    a[21] = 20'b00000000000000010101;
    a[22] = 20'b00000000000000010110;
    a[23] = 20'b00000000000000010111;
    a[24] = 20'b00000000000000011000;
    a[25] = 20'b00000000000000011001;
    a[26] = 20'b00000000000000011010;
    a[27] = 20'b00000000000000011011;
    a[28] = 20'b00000000000000011100;
    a[29] = 20'b00000000000000011101;
    a[30] = 20'b00000000000000011110;
    a[31] = 20'b00000000000000011111;
    a[32] = 20'b00000000000000100000;
    a[33] = 20'b00000000000000100001;
    a[34] = 20'b00000000000000100010;
    a[35] = 20'b00000000000000100011;
    a[36] = 20'b00000000000000100100;
    a[37] = 20'b00000000000000100101;
    a[38] = 20'b00000000000000100110;
    a[39] = 20'b00000000000000100111;
    a[40] = 20'b00000000000000101000;
    a[41] = 20'b00000000000000101001;
    a[42] = 20'b00000000000000101010;
    a[43] = 20'b00000000000000101011;
    a[44] = 20'b00000000000000101100;
    a[45] = 20'b00000000000000101101;
    a[46] = 20'b00000000000000101110;
    a[47] = 20'b00000000000000101111;
    a[48] = 20'b00000000000000110000;
    a[49] = 20'b00000000000000110001;
    a[50] = 20'b00000000000000110010;
    a[51] = 20'b00000000000000110011;
    a[52] = 20'b00000000000000110100;
    a[53] = 20'b00000000000000110101;
    a[54] = 20'b00000000000000110110;
    a[55] = 20'b00000000000000110111;
    a[56] = 20'b00000000000000111000;
    a[57] = 20'b00000000000000111001;
    a[58] = 20'b00000000000000111010;
    a[59] = 20'b00000000000000111011;
    a[60] = 20'b00000000000000111100;
    a[61] = 20'b00000000000000111101;
    a[62] = 20'b00000000000000111110;
    a[63] = 20'b00000000000000111111;

    C = 20'b00000000000000000000;

    R = 6'b000000;
    #10;

    R = 6'b000001;
    #10;
    
    R = 6'b100000;
    #10;

    R = 6'b110000;
    #10;

    R = 6'b111111;
    #10;

    $finish;

end

endmodule
